
---
"%test":
  ide-sidecar:
    connections:
      ccloud:
        control-plane-base-url: http://localhost:${quarkus.wiremock.devservices.port}
        id-token:
          exchange-uri: http://localhost:${quarkus.wiremock.devservices.port}/oauth/token
        control-plane-token:
          exchange-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/sessions
          check-jwt-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/check_jwt
        data-plane-token:
          exchange-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/access_tokens
        oauth:
          login-realm-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/login/realm
        resources:
          org-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/org/v2/organizations
          env-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/org/v2/environments
          lkc-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/cmk/v2/clusters?environment=%s
          sr-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/srcm/v3/clusters?environment=%s
          flink-compute-pools-uri: http://localhost:${quarkus.wiremock.devservices.port}/api/fcpm/v2/compute-pools?environment=%s
      confluent-local:
        resources:
          clusters-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/v3/clusters
          brokers-list-uri: http://localhost:${quarkus.wiremock.devservices.port}/v3/clusters/%s/brokers
          broker-adv-listeners-config-uri: http://localhost:${quarkus.wiremock.devservices.port}/v3/clusters/%s/brokers/%s/configs/advertised.listeners
          kafka-topic-uri: http://localhost:${quarkus.wiremock.devservices.port}/v3/clusters/%s/topics/%s
    grim-reaper:
      # Should we check for remaining living vs code processes at all, and exit() if none left?
      enabled: false
      # How often to check?
      interval-seconds: 60
    flink-language-service-proxy:
      url-pattern: ws://127.0.0.1:${quarkus.http.test-port}/fls-mock
    schema-fetch-error-ttl: 30
    schema-fetch-retry:
      max-retries: 3
    flink:
      url-pattern: http://localhost:${quarkus.wiremock.devservices.port}/flink.%s.%s.confluent.cloud
  quarkus:
    wiremock:
      devservices:
        enabled: true
    http:
      # 1 higher than the default port, to avoid conflicting with the main application.
      port: 26637
      test-port: 26637
    smallrye-openapi:
      # Unset the store-schema-directory to avoid storing
      # OpenAPI schemas with the test port.
      store-schema-directory: ""
    log:
      console:
        json: false

"%dev":
  ide-sidecar:
    access_token_filter:
      enabled: false
    grim-reaper:
      # Should we check for remaining living vs code processes at all, and exit() if none left?
      enabled: false
      # How often to check?
      interval-seconds: 60
  quarkus:
    log:
      console:
        json: false

vscode:
  extension:
    version: unknown
  version: unknown

ide-sidecar:
  api:
    group: gateway
    groupWithVersion: ${ide-sidecar.api.group}/${ide-sidecar.api.version}
    host: http://localhost:${quarkus.http.port}
    version: v1
  connections:
    ccloud:
      check-token-expiration:
        interval-seconds: 5
      control-plane-base-url: https://api.devel.cpdev.cloud
      control-plane-token:
        exchange-uri: https://api.devel.cpdev.cloud/sessions
        check-jwt-uri: https://api.devel.cpdev.cloud/check_jwt
        life-time-seconds: 300
      data-plane-token:
        exchange-uri: https://api.devel.cpdev.cloud/access_tokens
      id-token:
        exchange-uri: https://login.confluent-dev.io/oauth/token
        life-time-seconds: 60
      oauth:
        authorize-uri: https://login.confluent-dev.io/oauth/authorize
        client-id: cUmAgrkbAZSqSiy38JE7Ya3i7FwXmyUF
        login-realm-uri: https://api.devel.cpdev.cloud/login/realm
        redirect-uri: http://127.0.0.1:26636/gateway/v1/callback-vscode-docs
        # URI redirect to tell the VS Code extension if the auth flow completed successfully or not
        vscode-extension-uri: vscode://confluentinc.vscode-confluent/authCallback
        scope: email openid offline_access
      refresh-status-interval-seconds: 5
      refresh-token:
        absolute-lifetime-seconds: 28800
        max-refresh-attempts: 50
      resources:
        homepage-uri: https://devel.cpdev.cloud/
        org-list-uri: https://api.devel.cpdev.cloud/org/v2/organizations
        env-list-uri: https://api.devel.cpdev.cloud/org/v2/environments
        lkc-list-uri: https://api.devel.cpdev.cloud/cmk/v2/clusters?environment=%s
        sr-list-uri: https://api.devel.cpdev.cloud/srcm/v3/clusters?environment=%s
        flink-compute-pools-uri: https://api.devel.cpdev.cloud/fcpm/v2/compute-pools?environment=%s

    confluent-local:
      # We assume that the user is running the confluent-local image with
      # the configured defaults as follows.
      # https://github.com/confluentinc/kafka-images/blob/7.4.x/local/include/etc/confluent/docker/configureDefaults
      default:
        kafkarest-uri: http://localhost:8082
        kafkarest-hostname: rest-proxy
        cluster-name: confluent-local
        schema-registry-uri: http://localhost:8081
      refresh-status-interval-seconds: 5
      resources:
        clusters-list-uri: ${ide-sidecar.connections.confluent-local.default.kafkarest-uri}/v3/clusters
        brokers-list-uri: ${ide-sidecar.connections.confluent-local.default.kafkarest-uri}/v3/clusters/%s/brokers
        broker-adv-listeners-config-uri: ${ide-sidecar.connections.confluent-local.default.kafkarest-uri}/v3/clusters/%s/brokers/%s/configs/advertised.listeners
        kafka-topic-uri: ${outpost.connections.confluent-local.default.kafkarest-uri}/v3/clusters/%s/topics/%s

    direct:
      refresh-status-interval-seconds: 5
      timeout-seconds: 5
  flink:
    url-pattern: https://flink.%s.%s.confluent.cloud
  access_token_filter:
    excluded_paths:
      # Following needed by oauth
      - /api/login/realm
      - /gateway/v1/callback-vscode-docs
      - /
      # And finally, the handshake route itself.
      - /gateway/v1/handshake
  grim-reaper:
    # Should we check for remaining living vs code processes at all, and exit() if none left?
    enabled: true
    # How often to check?
    interval-seconds: 60
  flink-language-service-proxy:
    reconnect-attempts: 1
    url-pattern: wss://flinkpls.{{ region }}.{{ provider }}.devel.cpdev.cloud/lsp
  proxy:
    ccloud-api-control-plane-regex: "(/artifact.*)|(/fcpm/v2/compute-pools.*)|(/metadata/security/v2alpha1/authorize)"
    ccloud-api-flink-data-plane-regex: "(/sql/v1.*)"
  websockets:
    # How long do we allow a connection to be established w/o it saying HELLO?
    initial-grace-seconds: 60
    # ... and how often do we check?
    purge-interval-seconds: 60
  # Configuration set by the sidecar when instantiating the Kafka Admin client
  # (We may choose to allow connection-specific overrides in the future)
  admin-client-configs:
    "client.id": Confluent for VS Code sidecar ${vscode.extension.version} - Admin
    "default.api.timeout.ms": 5000
    "request.timeout.ms": 5000
  # Configuration set by the sidecar when instantiating the Kafka Consumer
  # (We may choose to allow connection-specific overrides in the future)
  consumer-client-configs:
    "client.id": Confluent for VS Code sidecar ${vscode.extension.version} - Consumer
    "session.timeout.ms": 45000
  # Configuration set by the sidecar when instantiating the Kafka Producer
  # (We may choose to allow connection-specific overrides in the future)
  producer-client-configs:
    acks: all
    "client.id": Confluent for VS Code sidecar ${vscode.extension.version} - Producer
  # Configuration set by the sidecar when instantiating Kafka record serializers and deserializers.
  # See https://github.com/confluentinc/schema-registry/blob/master/schema-serializer/src/main/java/io/confluent/kafka/serializers/AbstractKafkaSchemaSerDeConfig.java#L39
  # for a full list of available configs.
  serde-configs:
    # Use sidecar provided SR proxy as the schema registry URL
    # Should be unused by serializers since we pass the
    # SchemaRegistryClient instance to them directly.
    "schema.registry.url": ${ide-sidecar.api.host}
    # Disable auto-registering schemas, as we expect the schema to be registered
    # before the data is serialized.
    "auto.register.schemas": "false"
    # Do not try to fetch the latest version of the schema from the registry
    "use.latest.version": "false"
    "key.subject.name.strategy": "io.confluent.kafka.serializers.subject.TopicNameStrategy"
    "value.subject.name.strategy": "io.confluent.kafka.serializers.subject.TopicNameStrategy"
  cluster-proxy:
    # Exclude these HTTP headers when proxying requests to the remote cluster (Kafka or Schema Registry)
    # It shouldn't really hurt if we _don't_ exclude these headers, but it's just cleaner to do so.
    http-header-exclusions:
      - x-connection-id
      - x-cluster-id
      - x-ccloud-region
      - x-ccloud-provider
      - Authorization
      - Host
      - Connection
      # This may contradict UTF-8 decoding done in the proxy response processing
      # https://github.com/confluentinc/ide-sidecar/issues/102
      - Accept-Encoding
  webclient:
    connect-timeout-seconds: 10
  schema-fetch-error-ttl: 30
  schema-fetch-retry:
    initial-backoff-ms: 250
    max-backoff-ms: 5000
    timeout-ms: 10000
    max-retries: 5
  integration-tests:
    # cp-demo configs used by Confluent Platform integration tests
    cp-demo:
      tag: v7.7.1

quarkus:
  apicurio-registry:
    devservices:
      enabled: false
  application:
    name: ide-sidecar
  banner:
    enabled: false
  kafka:
    devservices:
      # We do not use the Quarkus Kafka devservices container to start the Kafka cluster
      enabled: false
  log:
    min-level: INFO
    category:
      "org.apache.kafka.clients":
        level: ERROR
      "org.apache.kafka.common":
        level: ERROR
      "io.confluent.kafka.serializers":
        level: ERROR
      "io.qua.hib.val.deployment":
        level: INFO
      "io.qua.dep.ste.ReflectiveHierarchyStep":
        level: INFO
  http:
    host: 127.0.0.1
    port: 26636
    cors:
      ~: true
      origins: https://login.confluent-dev.io,https://login-stag.confluent-dev.io,https://login.confluent.io
  jackson:
    fail-on-unknown-properties: true
  native:
    additional-build-args: --initialize-at-run-time=io.confluent.idesidecar.restapi.auth.CCloudOAuthConfig\,io.confluent.idesidecar.restapi.auth.CCloudOAuthContext\,io.confluent.ide.sidecar.restapi.util.WebClientFactory\,org.apache.kafka.common.security.authenticator.SaslClientAuthenticator\,org.apache.avro.file.DataFileWriter\,io.confluent.kafka.schemaregistry.avro.AvroSchemaUtils\,com.github.luben.zstd
    resources:
      includes: templates/callback.html,templates/callback_failure.html,templates/default.html,templates/reset_password.html,feature-flag-defaults.json
  smallrye-health:
    root-path: /gateway/v1/health
    openapi:
      included: true
  ssl:
    native: true
  smallrye-openapi:
    path: /openapi
    info-title: Confluent ide-sidecar API
    store-schema-directory: src/generated/resources/
    info-version: ${quarkus.application.version}
    info-description: API for the Confluent ide-sidecar, part of Confluent for VS Code
    info-terms-of-service: Your terms here
    info-contact-email: vscode@confluent.io
    info-contact-name: Confluent for VS Code Support
    info-contact-url: https://confluent.io/contact
  smallrye-graphql:
    print-data-fetcher-exception: true
    root-path: /gateway/v1/graphql
    show-runtime-exception-message:
      -  io.confluent.idesidecar.restapi.exceptions.ConnectionNotFoundException
      -  io.confluent.idesidecar.restapi.exceptions.ResourceFetchingException
  scheduler:
    start-mode: forced
  swagger-ui:
    # By default, enable the Swagger UI in dev and test modes, but not during normal package builds.
    path: /swagger-ui
    always-include: false
  vertx:
    # Disable file caching in Vert.X since the native executable includes the path of the tmp dir
    # of the machine where the native image was built.
    caching: false
  kerberos:
    devservices:
      enabled: false

# Hide the /internal/kafka route from the OpenAPI spec
mp:
  openapi:
    scan:
      exclude:
        classes: >
          io.confluent.idesidecar.restapi.kafkarest.ClusterV3ApiImpl,
          io.confluent.idesidecar.restapi.kafkarest.TopicConfigV3ApiImpl,
          io.confluent.idesidecar.restapi.kafkarest.PartitionV3ApiImpl,
          io.confluent.idesidecar.restapi.kafkarest.RecordsV3ApiImpl,
          io.confluent.idesidecar.restapi.kafkarest.TopicV3ApiImpl
